// do I need a reset? 

module t_flipflop (
    input D, CLK, T,

//should these be reg?
    output reg Q,
    output NotQ
);

//mux instance
// takes T as enable switch, Q and NotQ as inputs

//dflipflop instance


endmodule