module mux(

);

endmodule
