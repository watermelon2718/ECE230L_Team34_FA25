module top (
    input [15:0] sw,
    output [15:0] led
);
    wire muxOut;

    mux mux_inst (
        //assign stuff
    );

    demux demux_inst (
        //assign stuff
    );

endmodule
