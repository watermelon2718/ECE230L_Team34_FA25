module top(
    input btnU, btnC,
    output [6:0] led
);

//ripple counter and modulo divider inst here

endmodule