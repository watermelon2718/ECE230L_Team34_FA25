module d_latch(
    input D, E,
    output Q, NotQ
);

    // Will contain D-Latch behavior

endmodule

