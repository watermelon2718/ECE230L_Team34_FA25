module top (
    input sw[9:0],
    output led[13:0]
);



endmodule